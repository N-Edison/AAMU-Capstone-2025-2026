.title KiCad schematic
.include "/Users/nemo/Desktop/Capstone Project 2025-2026/BJT OP-AMP 2025-2026/"
.model Q1.BJT2N3904 NPN
.model Q2.BJT2N3904 NPN
.model Q9.BJT2N3904 NPN
.model Q7.BJT2N3906 PNP
.model Q3.BJT2N3904 NPN
.model Q5.BJT2N3904 NPN
.model Q4.BJT2N3906 PNP
.model Q8.BJT2N3906 PNP
.model Q6.BJT2N3904 NPN
.save all
.probe alli
.probe p(R13)
.probe p(R12)
.probe p(R2)
.probe p(R11)
.probe p(Q1)
.probe p(Q2)
.probe p(C1)
.probe p(XRV2)
.probe p(R9)
.probe p(R5)
.probe p(XRV3)
.probe p(R7)
.probe p(R8)
.probe p(Q9)
.probe p(R1)
.probe p(XRV1)
.probe p(Q7)
.probe p(R3)
.probe p(Q3)
.probe p(R4)
.probe p(Q5)
.probe p(R14)
.probe p(R6)
.probe p(C2)
.probe p(Q4)
.probe p(Q8)
.probe p(Q6)
R13 VDD Net-_Q4-E_ 10
R12 VDD Net-_Q7-E_ 10
R2 Net-_Q2-E_ VSS 10
R11 Net-_Q1-E_ VSS 10
Q1 Net-_D1-K_ Bias Net-_Q1-E_ Q1.BJT2N3904
Q2 Bias Bias Net-_Q2-E_ Q2.BJT2N3904
C1 Net-_C1-Pad1_ OUT 0.001u
XRV2 Net-_R9-Pad2_ Net-_Q5-C_ Net-_R8-Pad2_ potentiometer
R9 Net-_Q6-E_ Net-_R9-Pad2_ 100
R5 Net-_Q6-E_ Net-_Q5-C_ 220
XRV3 unconnected-_RV3-Pad1_ Net-_R14-Pad2_ Net-_C1-Pad1_ potentiometer
R7 Net-_Q9-E_ VSS 10
R8 Net-_Q3-E_ Net-_R8-Pad2_ 100
Q9 OUT Bias Net-_Q9-E_ Q9.BJT2N3904
R1 /TRIM Bias 680
XRV1 unconnected-_RV1-Pad1_ VDD /TRIM potentiometer
Q7 Net-_Q7-E_ /Mirror /Mirror Q7.BJT2N3906
R3 Net-_Q3-E_ Net-_Q5-C_ 220
Q3 /Mirror V- Net-_Q3-E_ Q3.BJT2N3904
R4 Net-_Q5-E_ VSS 10
Q5 Net-_Q5-C_ Bias Net-_Q5-E_ Q5.BJT2N3904
R14 /Difference Net-_R14-Pad2_ 10
R6 VDD Net-_Q8-E_ 10
C2 VDD VSS 10u
Q4 Net-_Q4-E_ /Mirror /Difference Q4.BJT2N3906
Q8 Net-_Q8-E_ /Difference OUT Q8.BJT2N3906
Q6 /Difference V+ Net-_Q6-E_ Q6.BJT2N3904
.end
